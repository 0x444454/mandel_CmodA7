// 256-entry palette: iter8 -> RGB888.
//
// Change colors here.
// NOTE: The first color is usually supposed to be Black (Mandelbrot proper set), but feel free to break the rules ;-)

module palette_rom_256x12(
    input  logic        clk,
    input  logic [7:0]  addr,
    output logic [23:0] rgb888
);

    // Synthesis hint: prefer BRAM for the palette.
    (* rom_style = "block" *) logic [23:0] rom [0:255];

    initial begin
        rom = '{
            24'h000000, 24'h001155, 24'h002288, 24'h113399, 24'h224488, 24'h445588, 24'h666677, 24'h888866, 24'hBBAA55, 24'hEEBB55, 24'hFFCC66, 24'hFFDD99, 24'hEEDDAA, 24'hEEDDBB, 24'hDDDDCC, 24'hDDDDDD,
            24'hDDCCDD, 24'hD7C1DD, 24'hD2B5DD, 24'hCCAADD, 24'hCC99DD, 24'hCC88DD, 24'hCC77DD, 24'hCC66DD, 24'hCC55DD, 24'hCC44DD, 24'hBB33CC, 24'hBB22CC, 24'hB51CCC, 24'hB017CC, 24'hAA16CC, 24'hA414CC,
            24'h9F12CC, 24'h9717D2, 24'h901DD7, 24'h8824D9, 24'h7F2CDB, 24'h7733DD, 24'h6C3EDD, 24'h604ADD, 24'h5555DD, 24'h5566EE, 24'h4A71EE, 24'h3E7DEE, 24'h3388EE, 24'h3399EE, 24'h2299EE, 24'h22AAEE,
            24'h22BBEE, 24'h22BBFF, 24'h22C4FF, 24'h22CCFF, 24'h22D4FF, 24'h22DDFF, 24'h2DE3FF, 24'h39E8FF, 24'h44EEFF, 24'h55EEFF, 24'h66EEFF, 24'h77F4FF, 24'h88F9FF, 24'h99FFFF, 24'hAAFFFF, 24'hBBFFFF,
            24'hC6FFFF, 24'hD2FFFF, 24'hD1FFFF, 24'hD0FFFF, 24'hCFFFFF, 24'hCEFFFF, 24'hCDFFFF, 24'hC7FFFF, 24'hC1FFFF, 24'hBBFFFF, 24'hAAFFFF, 24'h99FFFF, 24'h88FFFF, 24'h88EEFF, 24'h77EEFF, 24'h66EEFF,
            24'h55EEFF, 24'h4AEEFF, 24'h3EEEFF, 24'h3AE8F9, 24'h37E3F4, 24'h36E1EC, 24'h34DFE5, 24'h34DEDD, 24'h33DED4, 24'h39D8CC, 24'h3ED2C3, 24'h46D0BB, 24'h4DCEB2, 24'h55CCAA, 24'h55CC99, 24'h66CC99,
            24'h66BB88, 24'h77BB77, 24'h77BB66, 24'h88BB66, 24'h88BB55, 24'h99AA55, 24'h9FAA4A, 24'hA4AA3E, 24'hAAAA33, 24'hAAAA22, 24'hB0AA1C, 24'hB5AA17, 24'hBBAA11, 24'hCCAA11, 24'hD2AA0B, 24'hD7AA06,
            24'hDAAC05, 24'hDEAF04, 24'hE1B103, 24'hE4B403, 24'hE7B602, 24'hEBB901, 24'hECBD01, 24'hECC101, 24'hEDC400, 24'hEDC800, 24'hEDCD00, 24'hEED200, 24'hEED800, 24'hF2D900, 24'hF6DA00, 24'hFBDC00,
            24'hFCE200, 24'hFEE800, 24'hFEE700, 24'hFEE600, 24'hFEE500, 24'hFEE400, 24'hFEE300, 24'hFEE200, 24'hFFE200, 24'hFFE100, 24'hFFE000, 24'hFFDF00, 24'hFFDE00, 24'hFFD800, 24'hFFD200, 24'hFFCC00,
            24'hFFC100, 24'hFFB500, 24'hFFAA00, 24'hFF9900, 24'hFF8800, 24'hFF7D00, 24'hFF7100, 24'hFF6600, 24'hFF5B00, 24'hFF4F00, 24'hFF4600, 24'hFF3C00, 24'hFF3300, 24'hFF2B00, 24'hFF2200, 24'hFF1A00,
            24'hFF1100, 24'hFF0900, 24'hFC0700, 24'hF80500, 24'hF50400, 24'hF10200, 24'hED0203, 24'hE90107, 24'hE5010A, 24'hE1000E, 24'hDA000F, 24'hD30010, 24'hCB0010, 24'hC30011, 24'hBD0011, 24'hB60011,
            24'hB00011, 24'hAA0011, 24'hAA0022, 24'h9F0022, 24'h930022, 24'h8A0022, 24'h800022, 24'h7D0024, 24'h7A0026, 24'h760028, 24'h73002A, 24'h70002D, 24'h6C002F, 24'h690031, 24'h670031, 24'h650031,
            24'h620032, 24'h600032, 24'h5E0032, 24'h5C0032, 24'h590033, 24'h570033, 24'h550033, 24'h530033, 24'h510033, 24'h4F0033, 24'h4C0033, 24'h4A0033, 24'h480033, 24'h460033, 24'h440033, 24'h420233,
            24'h400433, 24'h3E0633, 24'h3C0833, 24'h3B0933, 24'h390B33, 24'h370D33, 24'h350F33, 24'h350F36, 24'h34103A, 24'h34103D, 24'h331141, 24'h301142, 24'h2D1142, 24'h2A1142, 24'h281143, 24'h251144,
            24'h231144, 24'h221144, 24'h201144, 24'h1E1144, 24'h1D1144, 24'h1B1144, 24'h191144, 24'h181144, 24'h161144, 24'h141144, 24'h131144, 24'h121144, 24'h101144, 24'h0F1144, 24'h0D1144, 24'h0C1144,
            24'h0A1144, 24'h091144, 24'h071144, 24'h061144, 24'h041144, 24'h031144, 24'h011144, 24'h001144, 24'h001144, 24'h001144, 24'h001144, 24'h001144, 24'h001144, 24'h001144, 24'h001144, 24'h001144
        };
    end

    always_ff @(posedge clk) begin
        rgb888 <= rom[addr];
    end

endmodule
